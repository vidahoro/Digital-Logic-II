library verilog;
use verilog.vl_types.all;
entity alu_test_vlg_vec_tst is
end alu_test_vlg_vec_tst;
