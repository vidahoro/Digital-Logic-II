library verilog;
use verilog.vl_types.all;
entity rom_128x8_sync_vlg_vec_tst is
end rom_128x8_sync_vlg_vec_tst;
