library verilog;
use verilog.vl_types.all;
entity rw_96x8_sync_vlg_vec_tst is
end rw_96x8_sync_vlg_vec_tst;
