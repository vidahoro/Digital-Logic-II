library verilog;
use verilog.vl_types.all;
entity rom_test_vlg_vec_tst is
end rom_test_vlg_vec_tst;
